`timescale 1ns / 1ps

// register file

module reg_file(
input clk,
input reset,
input write_en,
input [4:0] rd_addr1,
input [4:0] rd_addr2,
input [4:0] wr_addr,
input [31:0] wr_data,
output [31:0] rd_data1,
output [31:0] rd_data2
);

reg [31:0] reg_file [31:0];
integer k;
assign rd_data1=reg_file[rd_addr1];
assign rd_data2=reg_file[rd_addr2];
always @ (posedge clk)
begin 
     if (reset)
	  begin
//	       for(k=0;k<32;k=k+1)
            reg_file[0]= 32'b00000010001100101000000000100001;
				reg_file[1]= 32'b00000010001100101000000000100001;
				reg_file[2]= 32'b00000010001100101000000000100001;
				reg_file[3]= 32'b00000010001100101000000000100001;
				reg_file[4]= 32'b00000010001100101000000000100001;
				reg_file[5]= 32'b00000010001100101000000000100001;
				reg_file[6]= 32'b00000010001100101000000000100001;
				reg_file[7]= 32'b00000000000000000000000000001010;
				reg_file[8]= 32'b00000000000000000000000000001010;
				reg_file[9]= 32'b00000000000000000000000000001010;
				reg_file[10]= 32'b00000000000000000000000000001010;
				reg_file[11]= 32'b00000000000000000000000000001010;
				reg_file[12]= 32'b00000000000000000000000000001010;
				reg_file[13]= 32'b00000000000000000000000000001010;
				reg_file[14]= 32'b00000000000000000000000000001010;
				reg_file[15]= 32'b00000000000000000000000000001010;
				reg_file[16]= 32'b00000000000000000000000000001010;
				reg_file[17]= 32'b00000000000000000000000000001010;
				reg_file[18]= 32'b00000000000000000000000000001010;
				reg_file[19]= 32'b00000000000000000000000000001010;
				reg_file[20]= 32'b00000000000000000000000000001010;
				reg_file[21]= 32'b00000000000000000000000000001010;
				reg_file[22]= 32'b00000000000000000000000000001010;
				reg_file[23]= 32'b00000000000000000000000000001010;
				reg_file[24]= 32'b00000000000000000000000000001010;
				reg_file[25]= 32'b00000000000000000000000000001010;
				reg_file[26]= 32'b00000000000000000000000000001010;
				reg_file[27]= 32'b00000000000000000000000000001010;
				reg_file[28]= 32'b00000000000000000000000000001010;
				reg_file[29]= 32'b00000000000000000000000000001010;
				reg_file[30]= 32'b00000000000000000000000000001010;
				reg_file[31]= 32'b00000000000000000000000000001010;
			
	   end
	  else if(write_en)
	  reg_file[wr_addr]=wr_data;
end
endmodule

